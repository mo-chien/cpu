`timescale 1ns / 1ps
`include "ALU.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/04/21 09:44:22
// Design Name: 
// Module Name: ALU_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ALU_sim(

    );
    reg [31:0]    ALU_DA;
    reg [31:0]    ALU_DB;
    reg [3:0]     ALUCLT;
    wire          ALU_ZERO;
    wire          ALU_OverFlow;
    wire [31:0]   ALU_DC;
    ALU u_ALU(
        .ALU_DA       ( ALU_DA       ),
        .ALU_DB       ( ALU_DB       ),
        .ALUCLT       ( ALUCLT       ),
        .ALU_ZERO     ( ALU_ZERO     ),
        .ALU_OverFlow ( ALU_OverFlow ),
        .ALU_DC       ( ALU_DC       )
    );


    initial begin
        $dumpfile("ALU_wave.vcd");
        $dumpvars;
        ALU_DA=32'b0000_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0000_0000_0001_0001_0001_1111_0001_0000;
        ALUCLT=4'b0000;
        #10
        ALU_DA=32'b0000_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0000_0000_1110_1110_1110_0000_0000_0001;
        ALUCLT=4'b1000;
        #10

        ALU_DA=32'b0000_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0000_0000_0000_0000_0000_0000_0001_0000;
        ALUCLT=4'b0001;
        #10

        ALU_DA=32'b1011_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0100_1111_0011_0001_0001_1111_1110_1111;
        ALUCLT=4'b0010;
        #10
        ALU_DA=32'b0100_1111_0011_0001_0001_1111_1110_1111;
        ALU_DB=32'b1011_0000_1110_1110_1110_0000_0000_0001;
        ALUCLT=4'b0010;
        #10
        ALU_DA=32'b0100_1111_0011_0001_0001_1111_1110_1111;
        ALU_DB=32'b0000_0000_1110_1110_1110_0000_0000_0001;
        ALUCLT=4'b0010;
        #10 
        ALU_DA=32'b1000_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b1100_1111_0011_0001_0001_1111_1110_1111;
        ALUCLT=4'b0010;
        #10 

        ALU_DA=32'b0100_1111_0011_0001_0001_1111_1110_1111;
        ALU_DB=32'b1011_0000_1110_1110_1110_0000_0000_0001;
        ALUCLT=4'b0011;
        #10
        ALU_DA=32'b1011_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0100_1111_0011_0001_0001_1111_1110_1111;
        ALUCLT=4'b0011;
        #10 

        ALU_DA=32'b1011_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0100_1111_0011_0001_0001_1111_1110_1111;
        ALUCLT=4'b0100;
        #10

        ALU_DA=32'b0000_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0000_0000_0000_0000_0000_0000_0001_0000;
        ALUCLT=4'b0101;
        #10    
        ALU_DA=32'b1000_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0000_0000_0000_0000_0000_0000_0001_0000;
        ALUCLT=4'b0101;
        #10

        ALU_DA=32'b0000_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0000_0000_0000_0000_0000_0000_0001_0000;
        ALUCLT=4'b1101;
        #10    
        ALU_DA=32'b1000_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0000_0000_0000_0000_0000_0000_0001_0000;
        ALUCLT=4'b1101;
        #10

        ALU_DA=32'b1011_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0100_1111_0011_0001_0001_1111_1110_1111;
        ALUCLT=4'b0110;
        #10 

        ALU_DA=32'b1011_0000_1110_1110_1110_0000_0000_0001;
        ALU_DB=32'b0100_1111_0011_0001_0001_1111_1110_1111;
        ALUCLT=4'b0111;
        #10
        $finish;              
    end


endmodule

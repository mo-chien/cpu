module uart_tx (
    
);

endmodule //uart_tx